* analysis type *
.tran 1ns 100ns 0ns

* 
* input sources *
*V1 100 0 DC 5

*V2 200 0 PWL ( 0n 2.0 0.00000000005n 0 5n 0.0 5.00000000005n 2.0 10n 2.0 10.00000000005n 0.0 15n 0.0 15.00000000005n 2.0 20n 2 20.00000000005n 0.0 25n 0.0 25.00000000005n 2.0 30n 2.0 30.00000000005n 0.0 40n 0.0 40.00000000005n 2.0 50n 2.0 50.00000000005n 0.0 60n 0.0 60.00000000005n 2.0 70n 2.0 70.00000000005n 0.0 80n 0.0 80.00000000005n 2.0 90n 2.0 90.00000000005n 0.0 100n 0.0 100.00000000005n 2.0)

*V3 300 0 DC 0

V1 100 0 PULSE (2 0 0 .0000001ns 0.0000001ns 10ns 20ns)
V2 200 0 PULSE (0 2 0 .0000001ns 0.0000001ns 20ns 40ns)
V3 300 0 PULSE (2 0 0 .0000001ns 0.0000001ns 50ns 100ns)
* resistors to ground *
r1 100 0 1Meg
r2 200 0 1Meg
r3 300 0 1Meg

rload1 400 0 1Meg

*
* adc_bridge blocks *
aconverter1 [100 200 300]  [1 2 3] adc_bridge1

.model adc_bridge1 adc_bridge ( in_low =0.3 in_high =0.7
+ rise_delay =1.0e-12 fall_delay =1.0e-12)

a3 [1] [2] [3] [4] ff

a4 [4] [5] inv
.model ff flipflop(instance_id = 13 rise_delay = 1.0e-12 fall_delay = 1.0e-12 stop_time= 90.0e-9)
.model inv inverter(instance_id = 14 rise_delay = 1.0e-12 fall_delay = 1.0e-12 stop_time= 90.0e-9)
* dac_bridge blocks *
aconverter2 [4] [400] dac_bridge1

.model dac_bridge1 dac_bridge( out_low=0.25 out_high=5.0 
+out_undef=1.8 t_rise=0.5e-9 t_fall=0.5e-9) 

.end

