* analysis type *
.tran 1us 200us 0us

* 
* input sources *
*V1 100 0 PWL ( 0u 0 0.0000000005u 5.0 10u 5.0 10.00000000005u 0.0 20u 0.0 20.00000000005u 0.0 30u 0.0 30.00000000005u 0.0 40u 0.0 40.00000000005u 0.0 50u 0.0 50.00000000005u 0.0 60u 0.0 60.00000000005u 0.0 70u 0.0 70.00000000005u 0.0 80u 0.0 80.00000000005u 0.0 90u 0.0 90.00000000005u 0.0 100u 0.0)
*V1 100 0 DC 2.0
*V2 200 0 PWL ( 0u 2.0 0.00000000005u 0 5u 0.0 5.00000000005u 2.0 10u 2.0 10.00000000005u 0.0 15u 0.0 15.00000000005u 2.0 20u 2 20.00000000005u 0.0 25u 0.0 25.00000000005u 2.0 30u 2.0 30.00000000005u 0.0 40u 0.0 40.00000000005u 2.0 50u 2.0 50.00000000005u 0.0 60u 0.0 60.00000000005u 2.0 70u 2.0 70.00000000005u 0.0 80u 0.0 80.00000000005u 2.0 90u 2.0 90.00000000005u 0.0 100u 0.0 100.00000000005u 2.0)
V1 200 0 PULSE (2 0 0 .0000001ns 0.0000001ns 70us 140us)
V2 100 0 PULSE (2 0 0 .0000001ns 0.0000001ns 10us 20us)


* resistors to ground *
r1 100 0 1Meg
r2 200 0 1Meg

*rload1 300 0 1Meg
rload2 400 0 1Meg
rload3 500 0 1Meg
*rload4 600 0 1Meg

*
* adc_bridge blocks *
aconverter1 [100 200]  [1 2] adc_bridge1

.model adc_bridge1 adc_bridge ( in_low =0.3 in_high =0.7
+ rise_delay =1.0e-12 fall_delay =1.0e-12)

ac1 [1] [2] [3 4 5 6] count1
ac2 [3] [4] [34] and
ac3 [5] [6] [56] or
.model and and_nghdl(instance_id=11 rise_delay = 1.0e-7 fall_delay = 1.0e-7 stop_time= 190.0e-6) 
.model or or_nghdl(instance_id=12 rise_delay = 1.0e-7 fall_delay = 1.0e-7 stop_time= 190.0e-6)
.model count1 counter(instance_id=10 rise_delay = 1.0e-7 fall_delay = 1.0e-7 stop_time= 190.0e-6)

* dac_bridge blocks *
aconverter2 [34 56] [400 500] dac_bridge1

.model dac_bridge1 dac_bridge( out_low=0.25 out_high=5.0 
+out_undef=1.8 t_rise=0.5e-9 t_fall=0.5e-9) 

.end
